** Profile: "SCHEMATIC1-5"  [ E:\Code\Assignments\3rd Term\Electric Circuit Lab\Az 5\5\5-schematic1-5.sim ] 

** Creating circuit file "5-schematic1-5.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of e:\orCad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 400u 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\5-SCHEMATIC1.net" 


.END
