** Profile: "SCHEMATIC1-asd"  [ E:\CODE\Electric Circuit Lab\az1-SCHEMATIC1-asd.sim ] 

** Creating circuit file "az1-SCHEMATIC1-asd.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of e:\orCad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\az1-SCHEMATIC1.net" 


.END
