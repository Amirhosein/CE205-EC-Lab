** Profile: "SCHEMATIC1-4"  [ E:\Code\Assignments\3rd Term\Electric Circuit Lab\Az 5\4\4-schematic1-4.sim ] 

** Creating circuit file "4-schematic1-4.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of e:\orCad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 40m 0 40u 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\4-SCHEMATIC1.net" 


.END
