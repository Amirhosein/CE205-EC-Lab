** Profile: "SCHEMATIC1-3"  [ E:\Code\Assignments\3rd Term\Electrical Circuit Lab\Session 10\3\3-schematic1-3.sim ] 

** Creating circuit file "3-schematic1-3.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of e:\orCad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 100m 0 100u 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\3-SCHEMATIC1.net" 


.END
