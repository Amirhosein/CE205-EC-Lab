** Profile: "SCHEMATIC1-1"  [ E:\Code\Assignments\3rd Term\Electrical-Circuit-Lab-Fall400\Session 9\1\1-schematic1-1.sim ] 

** Creating circuit file "1-schematic1-1.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of e:\orCad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_V2 0 5 0.1 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\1-SCHEMATIC1.net" 


.END
