** Profile: "SCHEMATIC1-4"  [ E:\CODE\ASSIGNMENTS\3RD TERM\ELECTRICAL-CIRCUIT-LAB-FALL400\SESSION 7\4\4-SCHEMATIC1-4.sim ] 

** Creating circuit file "4-SCHEMATIC1-4.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of e:\orCad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 100 0.1 1000k
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\4-SCHEMATIC1.net" 


.END
