** Profile: "SCHEMATIC1-1"  [ E:\CODE\Electric Circuit Lab\Az 3\1\1-SCHEMATIC1-1.sim ] 

** Creating circuit file "1-SCHEMATIC1-1.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of e:\orCad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\1-SCHEMATIC1.net" 


.END
