** Profile: "SCHEMATIC1-2"  [ E:\Code\Assignments\3rd Term\Electrical Circuit Lab\Session 10\2\2-SCHEMATIC1-2.sim ] 

** Creating circuit file "2-SCHEMATIC1-2.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of e:\orCad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 3m 0 3u 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\2-SCHEMATIC1.net" 


.END
