** Profile: "SCHEMATIC1-3-2"  [ E:\Code\Assignments\3rd Term\Electrical Circuit Lab\Session 10\3\3-schematic1-3-2.sim ] 

** Creating circuit file "3-schematic1-3-2.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of e:\orCad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 1000 0.001 30k
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\3-SCHEMATIC1.net" 


.END
