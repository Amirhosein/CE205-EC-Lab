** Profile: "SCHEMATIC1-3"  [ E:\Code\Assignments\3rd Term\Electric Circuit Lab\Az 6\3\3-schematic1-3.sim ] 

** Creating circuit file "3-schematic1-3.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of e:\orCad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 0.06ms 0 
.STEP LIN PARAM r 1k 30k 5k 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\3-SCHEMATIC1.net" 


.END
