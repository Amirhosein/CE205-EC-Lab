** Profile: "SCHEMATIC1-1"  [ e:\code\assignments\3rd term\electric circuit lab\az 5\1\1-schematic1-1.sim ] 

** Creating circuit file "1-schematic1-1.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of e:\orCad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 60ms 0 200 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\1-SCHEMATIC1.net" 


.END
