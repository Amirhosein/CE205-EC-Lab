** Profile: "SCHEMATIC1-4"  [ E:\CODE\ASSIGNMENTS\3RD TERM\ELECTRICAL CIRCUIT LAB\SESSION 10\4\4-SCHEMATIC1-4.sim ] 

** Creating circuit file "4-SCHEMATIC1-4.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of e:\orCad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 60m 0 20u 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\4-SCHEMATIC1.net" 


.END
