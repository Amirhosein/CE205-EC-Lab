** Profile: "SCHEMATIC1-3"  [ E:\Code\Assignments\3rd Term\Electrical-Circuit-Lab-Fall400\Session 7\3\3-schematic1-3.sim ] 

** Creating circuit file "3-schematic1-3.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of e:\orCad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 100 0.1 1000k
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\3-SCHEMATIC1.net" 


.END
