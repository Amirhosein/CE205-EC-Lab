** Profile: "SCHEMATIC1-asd"  [ E:\CODE\ASSIGNMENTS\3RD TERM\ELECTRICAL CIRCUIT LAB\SESSION 10\4\asdasd-SCHEMATIC1-asd.sim ] 

** Creating circuit file "asdasd-SCHEMATIC1-asd.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of e:\orCad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 3m 0 1u 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\asdasd-SCHEMATIC1.net" 


.END
