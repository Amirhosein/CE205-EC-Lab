** Profile: "SCHEMATIC1-6"  [ E:\Code\Assignments\3rd Term\Electrical-Circuit-Lab-Fall400\Session 8\6\6-schematic1-6.sim ] 

** Creating circuit file "6-schematic1-6.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of e:\orCad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 3m 0 10u 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\6-SCHEMATIC1.net" 


.END
